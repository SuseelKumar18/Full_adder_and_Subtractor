// Full Subtractor in Verilog 
module full_subtractor ( 
    input  wire a, b, bin,       // Inputs 
    output wire diff, borrow     // Outputs 
); 
 
    // Logic equations 
    assign diff   = a ^ b ^ bin;                  // Difference 
    assign borrow = (~a & b) | (~(a ^ b) & bin);  // Borrow logic 
 
endmodule